FB2/DEFAULT    BIAS (VER. 22)   * RULES NPN:AE PNP:AE RP:AE
* INSPICE Version 7.4   Freitag, 28. Januar 2000   8:59:44
.TEMP 27
.OPT NUMDGT=8 RELTOL=0.001 ABSTOL=1PA VNTOL=1UV LIMPTS=0 ITL1=400
+ ITL2=60 ITL4=10 ITL5=0 CHGTOL=0.001PC PIVTOL=1E-13 PIVREL=2E-4 GMIN=1E-13
+ DIGFREQ=100G DIGDRVZ=100K
VCC VCC 0 5V AC 1
R01 IP1 0 100K
R02 IP4 0 100K
R03 IP5 0 100K
R04 VCC IN3 100K
R05 VCC IN31 100K
VSUB SUB 0 0V
.AC DEC 10 1HZ 100MEGHZ
Q201 202 202 203 0 N1
Q202 203 203 0 0 N1
Q203 206 202 207 0 N1
Q204 206 209 204 0 P1
Q205 206 215 205 0 N8
Q206 208 208 0 0 N4 0.750
Q207 209 209 210 0 P1
Q208 211 206 209 0 P1
Q209 211 215 207 0 N1
Q210 212 212 214 0 P1
Q211 212 211 213 0 N1
Q212 IP5 212 216 0 P1
Q213 IN3 215 207 0 N1
Q214 IP4 212 218 0 P1
Q215 IN31 211 219 0 N1
Q216 IP1 212 220 0 P1
Q217 221 221 VCC 0 P1
Q218 221 208 0 0 N2
Q219 0 215 222 0 S1
Q220 VH 221 VCC 0 P1
Q221 224 208 0 0 N1
Q222 VH VH 222 0 N1
Q223 222 222 223 0 N1
Q224 224 224 223 0 P1
Q225 VCC 222 VBG 0 N4
Q226 0 224 VBG 0 P4
D201 0 VCC DTISN1 36.000
D202 0 VBG DTISN1 36.000
R201 VCC 201 RPN 200K
R202 201 202 RPN 200K
R203 205 207 RP 2.6K
R204 VCC 204 RP 2.8K
R205 207 208 RP 17.5K
R206 VCC 210 RP 2.8K
R207 VCC 214 RP 2.8K
R208 213 215 RP 2.8K
R209 215 0 RP 60K
R210 VCC 216 RP 2.8K
R212 VCC 218 RP 2.8K
R213 219 215 RP 2.8K
R214 VCC 220 RP 2.8K
XC201 0 211 0 KNIN PARAMS:AREA=14K
.SUBCKT KNIN AL1 N SUB PARAMS:AREA=1
CNI AL1 NVS {0.55F*AREA}
DSUB SUB NVS DSEPI {AREA}
VSENSE1 NVS N
.ENDS
.OP
.PROBE/CSDF
.MODEL N1 NPN (IS=3.67E-17 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=6M ISE=6E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=280 IRB=30U RBM=35 RE=2.4 RC=413
+ XTB=.5 EG=1.186 XTI=3.2 CJE=137F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9
+ ITF=25M CJC=103F VJC=500M MJC=305M XCJC=222M TR=44N CJS=485F VJS=655M MJS=396M
+ FC=700M TRC1=3M)
.MODEL P1 LPNP (IS=3.83E-16 BF=2.50E+02 NF=1 VAF=1.00E+02 IKF=80U ISE=0.5F
+ NE=1.46 BR=37 NR=1 VAR=30 IKR=90U ISC=0 NC=1.47 RB=312 RE=40 RC=550 XTB=-400M
+ EG=1.186 XTI=10.7 CJE=44F VJE=580M MJE=270M TF=14N XTF=500M VTF=600M ITF=1U
+ CJC=434F VJC=590M MJC=375M XCJC=0 TR=42N FC=700M CJS=1P VJS=690M MJS=420M)
.MODEL N8 NPN (IS=2.94E-16 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=48M ISE=48E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=45 IRB=240U RBM=6 RE=.3 RC=137 XTB=.5
+ EG=1.186 XTI=3.2 CJE=1.1P VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9 ITF=200M
+ CJC=324F VJC=500M MJC=305M XCJC=222M TR=44N CJS=900F VJS=655M MJS=396M FC=700M
+ TRC1=3M)
.MODEL N4 NPN (IS=1.47E-16 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=24M ISE=24E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=90 IRB=120U RBM=11 RE=.6 RC=196 XTB=.5
+ EG=1.186 XTI=3.2 CJE=488F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9 ITF=100M
+ CJC=202F VJC=500M MJC=305M XCJC=222M TR=44N CJS=730F VJS=655M MJS=396M FC=700M
+ TRC1=3M)
.MODEL N2 NPN (IS=7.34E-17 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=12M ISE=12E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=140 IRB=60U RBM=18 RE=1.2 RC=258
+ XTB=.5 EG=1.186 XTI=3.2 CJE=274F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9
+ ITF=50M CJC=154F VJC=500M MJC=305M XCJC=222M TR=44N CJS=619F VJS=655M MJS=396M
+ FC=700M TRC1=3M)
.MODEL S1 PNP (IS=3.67E-16 BF=2.50E+02 NF=1 VAF=1.20E+02 IKF=40U ISE=2.3E-16
+ NE=1.45 BR=700M NR=1 VAR=25 IKR=200U ISC=8F NC=1.35 RB=100 RE=40 RC=60
+ XTB=-500M EG=1.186 XTI=2.7 CJE=50F VJE=900M MJE=330M TF=16N XTF=500M VTF=800M
+ CJC=328F VJC=630M MJC=410M XCJC=24M TR=1.6U FC=700M)
.MODEL P4 LPNP (IS=1.53E-15 BF=2.50E+02 NF=1 VAF=1.00E+02 IKF=320U ISE=2.0F
+ NE=1.46 BR=37 NR=1 VAR=30 IKR=360U ISC=0 NC=1.47 RB=160 RE=6.4 RC=335
+ XTB=-400M EG=1.186 XTI=10.7 CJE=184F VJE=580M MJE=270M TF=14N XTF=500M
+ VTF=600M ITF=4U CJC=725F VJC=590M MJC=375M XCJC=0 TR=42N FC=700M CJS=1.6P
+ VJS=690M MJS=420M)
.MODEL DTISN1 D (IS=5.13E-14 IKF=6M N=1.18 BV=6.2 NBV=.5 RS=40 EG=1.186
+ XTI=3.2 CJO=928F VJ=680M M=430M FC=700M TBV1=350U)
.MODEL RPN RES (R=1.00E+00 TC1=5.155M TC2=9.31U)
.MODEL RP RES (R=1.00E+00 TC1=1.938M TC2=6.263U)
.MODEL DSEPI D (IS=10.03E-20 EG=1.206 XTI=1.5 CJO=0.07F VJ=0.68 M=0.39 BV=60)
.END
