* Incremental Netlister - Release : 1.83.1.4
* Netlist Time: Jun 26 15:40:42 1997
* ViewList: UNIspice cmos.sch schematic gate.sch UNImacro extracted
*           symbolic
* StopList: UNIspice UNImacro

*--------------------------------------------------------------------
* Sub-Circuit Netlist:
* Block  : Transconduttore
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:46 1997
*--------------------------------------------------------------------
.SUBCKT SUB0 IN N0 OUT N1
VV5 NET15 0 3
VI3 NET7 0 2.4
II0 NET9 0 500u
II1 NET11 0 500u
II2 NET13 0 1m
QQ3 NET15 NET7 NET21 0 C41 1
QQ1 NET18 N0 NET11 0 C41 1
QQ0 NET21 IN NET9 0 C41 1
QQ4 NET15 NET7 NET18 0 C41 1
QQ5 N1 NET18 NET13 0 C41 1
QQ12 OUT NET21 NET13 0 C41 1
RREE NET9 NET11 20
RR10 N1 NET15 2.8K
RR11 OUT NET15 2.8K
.ENDS SUB0


*--------------------------------------------------------------------
* Sub-Circuit Netlist:
* Block  : Phase_Shifter
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:47 1997
*--------------------------------------------------------------------
.SUBCKT SUB1 IN N0 OUT N1
RR3 N1 OUT 2.5K
* Cell : Transconduttore (bench_gyr)
XI2  NET11 NET6 N1 OUT SUB0
* Cell : Transconduttore (bench_gyr)
XI1  OUT N1 NET11 NET6 SUB0
CC1 N1 N0 1.778p
CC1A OUT IN 1.778p
CCL NET11 NET6 8.887p
CC0 OUT N1 8p
.ENDS SUB1


*--------------------------------------------------------------------
* Main Circuit Netlist:
* Block  : Test_phs_shf
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:47 1997
*--------------------------------------------------------------------
VV1 NET7 0 5 AC 1 SIN 0 10m 102.6MEG 0 0
RR7 0 IN 1
RR3 0 OUT 1
EE8 IN 0 NET7 0 1
EE2 OUT 0 NET3 NET11 1
* Cell : Phase_Shifter (bench_gyr)
XI0  NET7 0 NET3 NET11 SUB1

.ac DEC 101 10k 1.00G
.tran 1.0e-9 100.0e-9 0 1.0e-9
.OP 

.probe

*---------------------------------------------------------------
* Spice Model : C41
*---------------------------------------------------------------
.model C41 
+ NPN
+ IS=2.27E-018 BF=1.00E+002 BR=1.00E+000 NF=1.00E+000
+ NR=1.00E+000 TF=6.00E-012 TR=1.00E-008 XTF=1.00E+001
+ VTF=1.50E+000 ITF=6.87E-003 PTF=3.75E+001 VAF=4.50E+001
+ VAR=3.00E+000 IKF=9.23E-003 IKR=1.16E-003 ISE=8.27E-017
+ NE=2.00E+000 ISC=4.47E-017 NC=1.50E+000 RE=1.34E+001
+ RB=2.00E+002 IRB=0.00E+000 RBM=3.49E+001 RC=2.22E+002
+ CJE=1.06E-014 VJE=1.05E+000 MJE=1.60E-001 CJC=1.03E-014
+ VJC=8.60E-001 MJC=3.40E-001 XCJC=1.80E-001 CJS=9.69E-015
+ VJS=8.20E-001 MJS=3.20E-001 EG=1.17E+000 XTB=1.70E+000
+ XTI=3.00E+000 KF=0.00E+000 AF=1.00E+000 FC=5.00E-001
*
