*BIQU.FILTER: DEVICEMODELL*
.WIDTH OUT=80
.SUBCKT UA741 2 3 6
* 2=-E , 3=+E , 6=A *
VEE 4 0 DC -15
VCC 7 0 DC 15
R1 1 4 1K
R2 15 4 50K
R3 5 4 1K
R4 17 4 5K
R5 18 16 39K
R6 22 23 4.5K
R7 20 23 7.5K
R8 21 4 50K
R9 19 4 50
R10 24 6 25
R11 6 25 50
C 22 14 30P
Q1 9 3 10 NPN
Q2 12 13 10 PNP
Q3 9 2 11 NPN
Q4 14 13 11 PNP
Q5 12 15 1 NPN
Q6 14 15 5 NPN
Q7 7 12 15 NPN
Q8 9 9 7 PNP
Q9 13 9 7 PNP
Q10 13 16 17 NPN
Q11 16 16 4 NPN
Q12 18 18 7 PNP
Q13 14 19 4 NPN
Q14 20 14 21 NPN
Q15 22 18 7 PNP
Q16 22 23 20 NPN
Q17 20 21 19 NPN
Q18 22 24 6 NPN
Q19 7 22 24 NPQ
Q20 4 20 25 PNQ
Q21 6 6 23 NPN
.MODEL NPN NPN BF=160 RB=100 CJS=2P
+TF=0.3N TR=6N CJE=3P CJC=2P VAF=100
.MODEL NPQ NPN BF=160 RB=100 CJS=2P
+TF=0.3N TR=6N CJE=3P CJC=2P VAF=100 IS=2P
.MODEL PNP PNP BF=20 RB=20 TF=1N TR=20N
+CJE=6P CJC=4P VAF=100
.MODEL PNQ PNP BF=20 RB=20 TF=1N TR=20N
+CJE=6P CJC=4P VAF=100 IS=2P
.ENDS UA741
XOP1 2 0 3 UA741
XOP2 4 0 5 UA741
XOP3 6 0 7 UA741
R1 1 2 10K
R2 2 3 100K
R3 3 4 10K
R4 4 5 10K
R5 5 6 10K
R6 2 7 10K
C1 2 3 0.016U
C2 6 7 0.016U
VE 1 0 AC 1
.OP
.AC DEC 101 1 10MEG
.probe/CSDF
.END
