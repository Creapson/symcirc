
* Block  : Transconduttore
.SUBCKT SUB0 IN N0 OUT N1
VV5 NET15 0 3
VI3 NET7 0 2.4
II0 NET9 0 500u
II1 NET11 0 500u
II2 NET13 0 1m
QQ3 NET15 NET7 NET21 0 C41 1
QQ1 NET18 N0 NET11 0 C41 1
QQ0 NET21 IN NET9 0 C41 1
QQ4 NET15 NET7 NET18 0 C41 1
QQ5 N1 NET18 NET13 0 C41 1
QQ12 OUT NET21 NET13 0 C41 1
RREE NET9 NET11 20
RR10 N1 NET15 2.8K
RR11 OUT NET15 2.8K
.ENDS SUB0

V1 1 2 AC 1
Voff 2 0 DC 1.5
X1 1 2 3 4 SUB0

.ac DEC 101 10k 1.00G
.OP

.probe

*---------------------------------------------------------------
* Spice Model : C41
*---------------------------------------------------------------
.model C41 
+ NPN
+ IS=2.27E-018 BF=1.00E+002 BR=1.00E+000 NF=1.00E+000
+ NR=1.00E+000 TF=6.00E-012 TR=1.00E-008 XTF=1.00E+001
+ VTF=1.50E+000 ITF=6.87E-003 PTF=3.75E+001 VAF=4.50E+001
+ VAR=3.00E+000 IKF=9.23E-003 IKR=1.16E-003 ISE=8.27E-017
+ NE=2.00E+000 ISC=4.47E-017 NC=1.50E+000 RE=1.34E+001
+ RB=2.00E+002 IRB=0.00E+000 RBM=3.49E+001 RC=2.22E+002
+ CJE=1.06E-014 VJE=1.05E+000 MJE=1.60E-001 CJC=1.03E-014
+ VJC=8.60E-001 MJC=3.40E-001 XCJC=1.80E-001 CJS=9.69E-015
+ VJS=8.20E-001 MJS=3.20E-001 EG=1.17E+000 XTB=1.70E+000
+ XTI=3.00E+000 KF=0.00E+000 AF=1.00E+000 FC=5.00E-001
*
* Frequenz-Spannungswandler
v0 1 0 sffm 0 200mv 1khz 5 100hz
vp 7 0 15v
vm 8 0 -15v
x1 1 2 3 7 8 macro741
x2 5 0 6 7 8 macro741
r0 1 0 100
r1 2 3 100k
r2 2 0 100
r3 5 6 1meg
c1 3 4 180pF ic=15V
c2 5 6 4.7nF ic=-5.2V
d1 4 0 diode
d2 5 4 diode
.model diode d (is=7nA n=2 rs=0.8)
* Teilschaltung OP741
.subckt macro741    2    3    6    7     4
*                   -in  +in  out   vp    vm
i0 7 1 1uA
vm1 9 4 0 
vm2 8 4 0
f1 7 5 vm1 1k
f2 5 4 vm2 1k
r1 7 5 10meg
r2 5 4 10meg
q1 9 2 1 nn1
q2 8 3 1 nn1
q3 4 5 6 nn2
q4 7 5 6 nn3
.model nn1 pnp (is=1p)
.model nn2 pnp (is=1p bf=1meg cjc=1nF mjc=0 re=100 nf=0.3)
.model nn3 npn (is=1p bf=1meg cjc=1nF mjc=0 re=100 nf=0.3)
.ends macro741
* End Teilschaltung OP741
.tran 40uS 20mS uic
.print tran v(1) v(3) v(6)
.options itl5=15000 limpts=501
.probe
FB2/DEFAULT    BIAS (VER. 22)   * RULES NPN:AE PNP:AE RP:AE
* INSPICE Version 7.4   Freitag, 28. Januar 2000   8:59:44
.TEMP 27
.OPT NUMDGT=8 RELTOL=0.001 ABSTOL=1PA VNTOL=1UV LIMPTS=0 ITL1=400
+ ITL2=60 ITL4=10 ITL5=0 CHGTOL=0.001PC PIVTOL=1E-13 PIVREL=2E-4 GMIN=1E-13
+ DIGFREQ=100G DIGDRVZ=100K
VCC VCC 0 5V AC 1
R01 IP1 0 100K
R02 IP4 0 100K
R03 IP5 0 100K
R04 VCC IN3 100K
R05 VCC IN31 100K
VSUB SUB 0 0V
.AC DEC 10 1HZ 100MEGHZ
Q201 202 202 203 0 N1
Q202 203 203 0 0 N1
Q203 206 202 207 0 N1
Q204 206 209 204 0 P1
Q205 206 215 205 0 N8
Q206 208 208 0 0 N4 0.750
Q207 209 209 210 0 P1
Q208 211 206 209 0 P1
Q209 211 215 207 0 N1
Q210 212 212 214 0 P1
Q211 212 211 213 0 N1
Q212 IP5 212 216 0 P1
Q213 IN3 215 207 0 N1
Q214 IP4 212 218 0 P1
Q215 IN31 211 219 0 N1
Q216 IP1 212 220 0 P1
Q217 221 221 VCC 0 P1
Q218 221 208 0 0 N2
Q219 0 215 222 0 S1
Q220 VH 221 VCC 0 P1
Q221 224 208 0 0 N1
Q222 VH VH 222 0 N1
Q223 222 222 223 0 N1
Q224 224 224 223 0 P1
Q225 VCC 222 VBG 0 N4
Q226 0 224 VBG 0 P4
D201 0 VCC DTISN1 36.000
D202 0 VBG DTISN1 36.000
R201 VCC 201 RPN 200K
R202 201 202 RPN 200K
R203 205 207 RP 2.6K
R204 VCC 204 RP 2.8K
R205 207 208 RP 17.5K
R206 VCC 210 RP 2.8K
R207 VCC 214 RP 2.8K
R208 213 215 RP 2.8K
R209 215 0 RP 60K
R210 VCC 216 RP 2.8K
R212 VCC 218 RP 2.8K
R213 219 215 RP 2.8K
R214 VCC 220 RP 2.8K
XC201 0 211 0 KNIN PARAMS:AREA=14K
.SUBCKT KNIN AL1 N SUB PARAMS:AREA=1
CNI AL1 NVS {0.55F*AREA}
DSUB SUB NVS DSEPI {AREA}
VSENSE1 NVS N
.ENDS
.OP
.PROBE/CSDF
.MODEL N1 NPN (IS=3.67E-17 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=6M ISE=6E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=280 IRB=30U RBM=35 RE=2.4 RC=413
+ XTB=.5 EG=1.186 XTI=3.2 CJE=137F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9
+ ITF=25M CJC=103F VJC=500M MJC=305M XCJC=222M TR=44N CJS=485F VJS=655M MJS=396M
+ FC=700M TRC1=3M)
.MODEL P1 LPNP (IS=3.83E-16 BF=2.50E+02 NF=1 VAF=1.00E+02 IKF=80U ISE=0.5F
+ NE=1.46 BR=37 NR=1 VAR=30 IKR=90U ISC=0 NC=1.47 RB=312 RE=40 RC=550 XTB=-400M
+ EG=1.186 XTI=10.7 CJE=44F VJE=580M MJE=270M TF=14N XTF=500M VTF=600M ITF=1U
+ CJC=434F VJC=590M MJC=375M XCJC=0 TR=42N FC=700M CJS=1P VJS=690M MJS=420M)
.MODEL N8 NPN (IS=2.94E-16 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=48M ISE=48E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=45 IRB=240U RBM=6 RE=.3 RC=137 XTB=.5
+ EG=1.186 XTI=3.2 CJE=1.1P VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9 ITF=200M
+ CJC=324F VJC=500M MJC=305M XCJC=222M TR=44N CJS=900F VJS=655M MJS=396M FC=700M
+ TRC1=3M)
.MODEL N4 NPN (IS=1.47E-16 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=24M ISE=24E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=90 IRB=120U RBM=11 RE=.6 RC=196 XTB=.5
+ EG=1.186 XTI=3.2 CJE=488F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9 ITF=100M
+ CJC=202F VJC=500M MJC=305M XCJC=222M TR=44N CJS=730F VJS=655M MJS=396M FC=700M
+ TRC1=3M)
.MODEL N2 NPN (IS=7.34E-17 BF=1.10E+02 NF=1 VAF=2.50E+02 IKF=12M ISE=12E-18
+ NE=1.18 BR=10 NR=1 VAR=30 ISC=0 NC=2 RB=140 IRB=60U RBM=18 RE=1.2 RC=258
+ XTB=.5 EG=1.186 XTI=3.2 CJE=274F VJE=755M MJE=340M TF=440P XTF=38 VTF=2.9
+ ITF=50M CJC=154F VJC=500M MJC=305M XCJC=222M TR=44N CJS=619F VJS=655M MJS=396M
+ FC=700M TRC1=3M)
.MODEL S1 PNP (IS=3.67E-16 BF=2.50E+02 NF=1 VAF=1.20E+02 IKF=40U ISE=2.3E-16
+ NE=1.45 BR=700M NR=1 VAR=25 IKR=200U ISC=8F NC=1.35 RB=100 RE=40 RC=60
+ XTB=-500M EG=1.186 XTI=2.7 CJE=50F VJE=900M MJE=330M TF=16N XTF=500M VTF=800M
+ CJC=328F VJC=630M MJC=410M XCJC=24M TR=1.6U FC=700M)
.MODEL P4 LPNP (IS=1.53E-15 BF=2.50E+02 NF=1 VAF=1.00E+02 IKF=320U ISE=2.0F
+ NE=1.46 BR=37 NR=1 VAR=30 IKR=360U ISC=0 NC=1.47 RB=160 RE=6.4 RC=335
+ XTB=-400M EG=1.186 XTI=10.7 CJE=184F VJE=580M MJE=270M TF=14N XTF=500M
+ VTF=600M ITF=4U CJC=725F VJC=590M MJC=375M XCJC=0 TR=42N FC=700M CJS=1.6P
+ VJS=690M MJS=420M)
.MODEL DTISN1 D (IS=5.13E-14 IKF=6M N=1.18 BV=6.2 NBV=.5 RS=40 EG=1.186
+ XTI=3.2 CJO=928F VJ=680M M=430M FC=700M TBV1=350U)
.MODEL RPN RES (R=1.00E+00 TC1=5.155M TC2=9.31U)
.MODEL RP RES (R=1.00E+00 TC1=1.938M TC2=6.263U)
.MODEL DSEPI D (IS=10.03E-20 EG=1.206 XTI=1.5 CJO=0.07F VJ=0.68 M=0.39 BV=60)
.END.ende
* Incremental Netlister - Release : 1.83.1.4
* Netlist Time: Jun 26 15:40:42 1997
* ViewList: UNIspice cmos.sch schematic gate.sch UNImacro extracted
*           symbolic
* StopList: UNIspice UNImacro

*--------------------------------------------------------------------
* Sub-Circuit Netlist:
* Block  : Transconduttore
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:46 1997
*--------------------------------------------------------------------
.SUBCKT SUB0 IN N0 OUT N1
VV5 NET15 0 3
VI3 NET7 0 2.4
II0 NET9 0 500u
II1 NET11 0 500u
II2 NET13 0 1m
QQ3 NET15 NET7 NET21 0 C41 1
QQ1 NET18 N0 NET11 0 C41 1
QQ0 NET21 IN NET9 0 C41 1
QQ4 NET15 NET7 NET18 0 C41 1
QQ5 N1 NET18 NET13 0 C41 1
QQ12 OUT NET21 NET13 0 C41 1
RREE NET9 NET11 20
RR10 N1 NET15 2.8K
RR11 OUT NET15 2.8K
.ENDS SUB0


*--------------------------------------------------------------------
* Sub-Circuit Netlist:
* Block  : Phase_Shifter
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:47 1997
*--------------------------------------------------------------------
.SUBCKT SUB1 IN N0 OUT N1
RR3 N1 OUT 2.5K
* Cell : Transconduttore (bench_gyr)
XI2  NET11 NET6 N1 OUT SUB0
* Cell : Transconduttore (bench_gyr)
XI1  OUT N1 NET11 NET6 SUB0
CC1 N1 N0 1.778p
CC1A OUT IN 1.778p
CCL NET11 NET6 8.887p
CC0 OUT N1 8p
.ENDS SUB1


*--------------------------------------------------------------------
* Main Circuit Netlist:
* Block  : Test_phs_shf
* Library: bench_gyr
* Last Time Saved: Jun 26 15:39:47 1997
*--------------------------------------------------------------------
VV1 NET7 0 5 AC 1 SIN 0 10m 102.6MEG 0 0
RR7 0 IN 1
RR3 0 OUT 1
EE8 IN 0 NET7 0 1
EE2 OUT 0 NET3 NET11 1
* Cell : Phase_Shifter (bench_gyr)
XI0  NET7 0 NET3 NET11 SUB1

.ac DEC 101 10k 1.00G
.tran 1.0e-9 100.0e-9 0 1.0e-9
.OP 

.probe

*---------------------------------------------------------------
* Spice Model : C41
*---------------------------------------------------------------
.model C41 
+ NPN
+ IS=2.27E-018 BF=1.00E+002 BR=1.00E+000 NF=1.00E+000
+ NR=1.00E+000 TF=6.00E-012 TR=1.00E-008 XTF=1.00E+001
+ VTF=1.50E+000 ITF=6.87E-003 PTF=3.75E+001 VAF=4.50E+001
+ VAR=3.00E+000 IKF=9.23E-003 IKR=1.16E-003 ISE=8.27E-017
+ NE=2.00E+000 ISC=4.47E-017 NC=1.50E+000 RE=1.34E+001
+ RB=2.00E+002 IRB=0.00E+000 RBM=3.49E+001 RC=2.22E+002
+ CJE=1.06E-014 VJE=1.05E+000 MJE=1.60E-001 CJC=1.03E-014
+ VJC=8.60E-001 MJC=3.40E-001 XCJC=1.80E-001 CJS=9.69E-015
+ VJS=8.20E-001 MJS=3.20E-001 EG=1.17E+000 XTB=1.70E+000
+ XTI=3.00E+000 KF=0.00E+000 AF=1.00E+000 FC=5.00E-001
*
